/*=============================================================================
 * Title        : Moving average testbench
 *
 * File Name    : MOVING_AVE.sv
 * Project      : 
 * Designer     : toms74209200 <https://github.com/toms74209200>
 * Created      : 2023/05/05
 * License      : MIT License.
                  http://opensource.org/licenses/mit-license.php
 *============================================================================*/

`timescale 1ns/1ns

`define Comment(sentence) \
$display("%0s(%0d) %0s.", `__FILE__, `__LINE__, sentence)
`define MessageOK(name, value) \
$display("%0s(%0d) OK:Assertion %0s = %0d.", `__FILE__, `__LINE__, name, value)
`define MessageERROR(name, variable, value) \
$error("%0s(%0d) ERROR:Assertion %0s = %0d failed. %0s = %0d", `__FILE__, `__LINE__, name, value, name, variable)
`define ChkValue(name, variable, value) \
    if ((variable)===(value)) \
        `MessageOK(name, value); \
    else \
        `MessageERROR(name, variable, value);

module TB_MOVING_AVE ;

// Simulation module signal
bit         RESET_n;            //(n) Reset
bit         CLK;                //(p) Clock
bit         ASI_READY;          //(p) Avalon-ST sink data ready
bit         ASI_VALID = 0;      //(p) Avalon-ST sink data valid
bit [15:0]  ASI_DATA  = 0;      //(p) Avalon-ST sink data
bit         ASO_VALID;          //(p) Avalon-ST source data valid
bit [15:0]  ASO_DATA;           //(p) Avalon-ST source data
bit         ASO_ERROR;          //(p) Avalon-ST source error

// Parameter
parameter ClkCyc    = 10;       // Signal change interval(10ns/50MHz)
parameter ResetTime = 20;       // Reset hold time

// Data rom
bit [15:0] raw_data_rom[0:1023] = {
    16'h30F4,
    16'h3AAD,
    16'h8581,
    16'h637C,
    16'h58F1,
    16'h9135,
    16'h9F9A,
    16'h0269,
    16'h7211,
    16'hA559,
    16'h681B,
    16'h8C8A,
    16'hB6E9,
    16'h40F6,
    16'h3FF3,
    16'hDC75,
    16'h8B34,
    16'h93C9,
    16'hEA0A,
    16'hD238,
    16'h4523,
    16'hBC33,
    16'hA9D0,
    16'hD683,
    16'h2105,
    16'h9921,
    16'hFE04,
    16'h3518,
    16'hC489,
    16'h1025,
    16'hA9C3,
    16'h0773,
    16'h013F,
    16'h8AD2,
    16'h6905,
    16'h0AC8,
    16'h7EF7,
    16'h6E0D,
    16'h97CC,
    16'h608A,
    16'h176E,
    16'h4A2A,
    16'hA9E0,
    16'h1866,
    16'h40F8,
    16'h388A,
    16'hC074,
    16'hB968,
    16'hB04E,
    16'h2B0F,
    16'hA4DA,
    16'h0F5A,
    16'h7DB2,
    16'h7A1E,
    16'h144E,
    16'h7437,
    16'h05CA,
    16'h0EE1,
    16'h031F,
    16'hC33B,
    16'h091E,
    16'h5769,
    16'h4C27,
    16'h67AD,
    16'hC95E,
    16'hCD38,
    16'h7B21,
    16'h2CE9,
    16'h359D,
    16'hEFA2,
    16'hDE19,
    16'h2BCF,
    16'hC478,
    16'hD4C4,
    16'h60FA,
    16'h0A20,
    16'h6DD0,
    16'h99EF,
    16'hAE71,
    16'h8353,
    16'hB148,
    16'h6604,
    16'h5200,
    16'h1749,
    16'h9CE5,
    16'h923C,
    16'h662D,
    16'h1336,
    16'h6928,
    16'hBA71,
    16'hCB68,
    16'h5511,
    16'hE462,
    16'hC96E,
    16'h0473,
    16'hD5EB,
    16'hDBB5,
    16'h77CB,
    16'hD476,
    16'h8C1B,
    16'hCCC4,
    16'h6456,
    16'h7C89,
    16'h6D2D,
    16'h035D,
    16'h7CD7,
    16'h05DE,
    16'h5EA9,
    16'h0118,
    16'hC759,
    16'h3B65,
    16'h0F1C,
    16'hEE10,
    16'h939C,
    16'h5118,
    16'hA15C,
    16'h2140,
    16'h01A4,
    16'h7C7B,
    16'hF737,
    16'h739D,
    16'h3DE6,
    16'h5CD2,
    16'h8E72,
    16'h5848,
    16'h72B7,
    16'h20CB,
    16'hF515,
    16'h5326,
    16'h3525,
    16'hBF49,
    16'h3A17,
    16'h61DD,
    16'h1BD7,
    16'h352F,
    16'hDB81,
    16'h1F53,
    16'hDE0F,
    16'h995F,
    16'h7783,
    16'hD5B3,
    16'hA443,
    16'h6402,
    16'h4027,
    16'h6340,
    16'h4E70,
    16'hF5B1,
    16'h0EF3,
    16'h7430,
    16'h5FE5,
    16'h47DC,
    16'h743C,
    16'hE71A,
    16'h7B1E,
    16'h2293,
    16'h15E9,
    16'hC996,
    16'h2EC9,
    16'hF0FC,
    16'h2B04,
    16'hB94B,
    16'h77B9,
    16'h8FB5,
    16'h05CB,
    16'h4268,
    16'hD3A5,
    16'hD785,
    16'h0168,
    16'h0FCA,
    16'h4379,
    16'h065F,
    16'hE4AC,
    16'h3B20,
    16'hE3CB,
    16'hB97E,
    16'hF246,
    16'h0781,
    16'hE2B0,
    16'hD15D,
    16'hE0BF,
    16'h34E6,
    16'hD089,
    16'h83B3,
    16'hDF57,
    16'hD09A,
    16'h7EA1,
    16'hCF83,
    16'h7498,
    16'hB97E,
    16'h96A9,
    16'h46D6,
    16'hDD31,
    16'h5537,
    16'hA3A8,
    16'hF708,
    16'hCD24,
    16'hD967,
    16'h11C4,
    16'h848B,
    16'hBAB9,
    16'h1EA9,
    16'h17B1,
    16'hEF4C,
    16'h3CF3,
    16'hAE13,
    16'h8BCA,
    16'h8273,
    16'hEAC5,
    16'hB49D,
    16'hB893,
    16'h3FAD,
    16'h242A,
    16'h9819,
    16'h4DB5,
    16'hF3EB,
    16'h0B55,
    16'h4548,
    16'h7991,
    16'h3662,
    16'h63F4,
    16'h96D7,
    16'hC145,
    16'hA5E6,
    16'h67D9,
    16'h3CB5,
    16'h884E,
    16'hA823,
    16'h55B2,
    16'hA646,
    16'h3101,
    16'hAED5,
    16'hCDBC,
    16'hE318,
    16'hD3EA,
    16'hF0F8,
    16'hED62,
    16'hD3DD,
    16'hAC85,
    16'h6BB0,
    16'h7D7D,
    16'h7CF7,
    16'h8487,
    16'hD720,
    16'hC683,
    16'h6B7A,
    16'hC2B7,
    16'hD5BA,
    16'h8C66,
    16'h0325,
    16'h6882,
    16'hAB5F,
    16'hCAEC,
    16'hBB5C,
    16'h95D0,
    16'h764A,
    16'hADF6,
    16'h6D7F,
    16'hA8FD,
    16'h1BEC,
    16'hD9A1,
    16'h33DB,
    16'h07B5,
    16'h727B,
    16'hAFFB,
    16'h5559,
    16'h8E25,
    16'hBBCD,
    16'h03BA,
    16'h9991,
    16'h817B,
    16'h86F2,
    16'h6C3B,
    16'hF3BE,
    16'h1377,
    16'h8B1C,
    16'h1D4E,
    16'hBAFE,
    16'hE9C1,
    16'h4A2B,
    16'hEB00,
    16'h4D9B,
    16'h3109,
    16'h7723,
    16'h672B,
    16'hC1A1,
    16'h41D9,
    16'hF8CF,
    16'h343B,
    16'h621A,
    16'h11A2,
    16'h781F,
    16'h2AD2,
    16'h7B17,
    16'hFC2E,
    16'h6915,
    16'h4AC4,
    16'h22CA,
    16'hC188,
    16'h040A,
    16'hA426,
    16'h84C1,
    16'h5790,
    16'hC472,
    16'hBC07,
    16'h1813,
    16'hC7CA,
    16'hBB50,
    16'hA425,
    16'hFFF5,
    16'hA6B8,
    16'h4EAB,
    16'hC0CB,
    16'h17EB,
    16'h62F8,
    16'hB64E,
    16'h9C4F,
    16'h6F1B,
    16'h6903,
    16'h99B0,
    16'h61CF,
    16'h7ED0,
    16'h531D,
    16'h686B,
    16'h6393,
    16'h290B,
    16'hA836,
    16'h8F0E,
    16'h2C22,
    16'h3B21,
    16'hC330,
    16'h895D,
    16'h3ACC,
    16'h92B6,
    16'hE422,
    16'h2478,
    16'h7D17,
    16'h6B69,
    16'h2BB1,
    16'h4B31,
    16'h9A39,
    16'h965B,
    16'hE598,
    16'hE77D,
    16'h731C,
    16'h4D25,
    16'hD79A,
    16'hF223,
    16'h4B1B,
    16'h2865,
    16'h8CE3,
    16'h421E,
    16'h759E,
    16'hFBA2,
    16'h87BB,
    16'hF548,
    16'h10AD,
    16'hB5CA,
    16'h0C99,
    16'hD17D,
    16'h23D2,
    16'h36A2,
    16'hF8FC,
    16'h66B4,
    16'hBDE5,
    16'h4962,
    16'hDCAB,
    16'hF472,
    16'h475B,
    16'hD059,
    16'h6F2C,
    16'h3FF8,
    16'h9963,
    16'h1E77,
    16'hF74E,
    16'h9868,
    16'hC06F,
    16'hE089,
    16'h74AC,
    16'hB547,
    16'hCDA3,
    16'h763F,
    16'h510F,
    16'hC684,
    16'h7662,
    16'h96A1,
    16'hAFEB,
    16'hEA9D,
    16'h39BE,
    16'h009B,
    16'h95C9,
    16'h4CA2,
    16'hB21A,
    16'h3762,
    16'hEF31,
    16'h5AE5,
    16'h5794,
    16'hF258,
    16'h8468,
    16'h3D19,
    16'hB62E,
    16'h9E43,
    16'h969E,
    16'hB107,
    16'h5995,
    16'h57C9,
    16'hDEEE,
    16'hCA6E,
    16'hD882,
    16'hB335,
    16'h6BFF,
    16'hD14D,
    16'h8510,
    16'h37F8,
    16'h0051,
    16'h72BD,
    16'hDDFD,
    16'h3270,
    16'h882F,
    16'h1C3A,
    16'h6E89,
    16'hA5CA,
    16'hA6B5,
    16'h4630,
    16'h54CC,
    16'hC442,
    16'h5DAA,
    16'h95D4,
    16'hD531,
    16'h5B2D,
    16'h6B28,
    16'h789D,
    16'h0F5B,
    16'hD6EF,
    16'h839F,
    16'h21B3,
    16'h17A6,
    16'hE98F,
    16'h629A,
    16'h4554,
    16'h6883,
    16'hE77D,
    16'h9DD2,
    16'h670D,
    16'hB297,
    16'h29A6,
    16'hEDA5,
    16'hBC5D,
    16'h664B,
    16'h151F,
    16'hB1B8,
    16'hB58B,
    16'h22B1,
    16'hD24F,
    16'hA6E0,
    16'h5AC6,
    16'h4FAE,
    16'h41A7,
    16'h9861,
    16'h8D53,
    16'h934D,
    16'h425A,
    16'h2EA3,
    16'hE3D5,
    16'h4026,
    16'h67CC,
    16'hE93C,
    16'h86D0,
    16'h7A20,
    16'hF09E,
    16'h5CD4,
    16'hA080,
    16'hAE68,
    16'hDB7D,
    16'hCCD4,
    16'h0AD3,
    16'h6F63,
    16'hBB0D,
    16'h500A,
    16'hBCA7,
    16'h554D,
    16'hFA7E,
    16'hD35A,
    16'h1DE7,
    16'hF0FB,
    16'hE60E,
    16'h35C2,
    16'h5804,
    16'h990D,
    16'h6AFE,
    16'hBEE7,
    16'hBE94,
    16'hFE4C,
    16'h6010,
    16'hC7D1,
    16'h32F6,
    16'h14D6,
    16'hE4C0,
    16'hE41B,
    16'h1E2E,
    16'h18C6,
    16'hBFC4,
    16'hD4E1,
    16'hE91A,
    16'h6ECB,
    16'h38A7,
    16'h9519,
    16'h8F97,
    16'h51AC,
    16'h0944,
    16'h76B7,
    16'h21EB,
    16'h1846,
    16'h8D05,
    16'hB7B8,
    16'h1A46,
    16'h48F4,
    16'h057F,
    16'h1AE5,
    16'h08FB,
    16'h39BB,
    16'hB3EB,
    16'h4E7F,
    16'h58B8,
    16'hCD7C,
    16'h9BAF,
    16'hA7DB,
    16'hA517,
    16'hB98A,
    16'hB6DF,
    16'hDE6D,
    16'h3FDE,
    16'hA424,
    16'hB6E4,
    16'h01E6,
    16'h849F,
    16'h60D2,
    16'hBF5D,
    16'h250E,
    16'h4412,
    16'hBE8F,
    16'h14ED,
    16'h5865,
    16'hAA93,
    16'hE3C4,
    16'h9E1B,
    16'hE38E,
    16'hFE3A,
    16'h6701,
    16'hE18D,
    16'h05C4,
    16'hDA2C,
    16'hCEC5,
    16'h753E,
    16'hAD56,
    16'hD2A1,
    16'hA0DF,
    16'hB58D,
    16'hFABE,
    16'hEF71,
    16'hF4E7,
    16'h2D03,
    16'h044F,
    16'h58A8,
    16'hDFAF,
    16'hFBD0,
    16'h4B95,
    16'h063D,
    16'hE6E9,
    16'hE937,
    16'h2F99,
    16'h9FCE,
    16'h37DA,
    16'hE467,
    16'hF6B5,
    16'hB92D,
    16'hEC1C,
    16'h9A52,
    16'hA85F,
    16'h6B0C,
    16'hE486,
    16'h1139,
    16'hE283,
    16'hC042,
    16'h22C3,
    16'h4083,
    16'h5FF6,
    16'h8014,
    16'hBD18,
    16'h350F,
    16'hFE42,
    16'h2F20,
    16'hE354,
    16'h0657,
    16'hB4C1,
    16'hEA1B,
    16'hA9D9,
    16'hA74B,
    16'hE26F,
    16'hB584,
    16'h7A25,
    16'h0946,
    16'hA006,
    16'h8A3B,
    16'h7BC4,
    16'hBA05,
    16'h7C4B,
    16'h480D,
    16'h7EC8,
    16'hBBBF,
    16'h79D9,
    16'hC5A3,
    16'h1615,
    16'h0619,
    16'h1999,
    16'h6BC1,
    16'h107A,
    16'h4D84,
    16'hD09E,
    16'h4442,
    16'h7D51,
    16'hD2A9,
    16'h4F36,
    16'h2002,
    16'h859D,
    16'hD0E8,
    16'h1E16,
    16'h2207,
    16'h0B4E,
    16'hD911,
    16'h96E7,
    16'h2893,
    16'h664D,
    16'hD64A,
    16'h48AA,
    16'hCA0F,
    16'h8E9F,
    16'h7740,
    16'hE464,
    16'h248B,
    16'hBB59,
    16'h4CAC,
    16'hDCA4,
    16'h25EF,
    16'h5331,
    16'hD903,
    16'h9198,
    16'hCCF6,
    16'hE0DD,
    16'h5E5B,
    16'h65AE,
    16'h92FB,
    16'h8180,
    16'hBB23,
    16'h5357,
    16'hE92D,
    16'hD74F,
    16'h2611,
    16'hEB06,
    16'hE33D,
    16'h7CC2,
    16'h91FA,
    16'h9ED4,
    16'h7D72,
    16'hBB9E,
    16'h4FBF,
    16'h2782,
    16'h2E49,
    16'h5018,
    16'h6AEC,
    16'h4B18,
    16'hC8D6,
    16'h5599,
    16'h6802,
    16'hF185,
    16'h8FA8,
    16'h5064,
    16'hF3FC,
    16'h45BB,
    16'h104D,
    16'hDDAE,
    16'hFBF1,
    16'hEBB9,
    16'hABD8,
    16'h0EC4,
    16'h0708,
    16'h47F8,
    16'h5119,
    16'h7F2C,
    16'hDDCA,
    16'h9D5E,
    16'h98A8,
    16'h453C,
    16'hE2DF,
    16'h8E91,
    16'h65F2,
    16'h7394,
    16'h1D24,
    16'hE23E,
    16'hF7C0,
    16'hF35D,
    16'h90A7,
    16'hE85C,
    16'h6207,
    16'h2F0E,
    16'h9979,
    16'hFC44,
    16'h27C5,
    16'hD20C,
    16'h132B,
    16'h1763,
    16'hAD89,
    16'h8055,
    16'hB7FA,
    16'h5C49,
    16'h17E5,
    16'h7E10,
    16'h2E08,
    16'h781C,
    16'h39A9,
    16'h015B,
    16'h2142,
    16'h84CE,
    16'h13A0,
    16'hFDBC,
    16'hA2F2,
    16'hAB70,
    16'h0B7E,
    16'h55C4,
    16'h84AB,
    16'hB5E7,
    16'h3BD3,
    16'h980D,
    16'hDE51,
    16'h6317,
    16'hE10A,
    16'h16FA,
    16'h328D,
    16'h9F33,
    16'h3D67,
    16'h6505,
    16'hE41D,
    16'hA5DB,
    16'h4096,
    16'h31C7,
    16'hBB49,
    16'hFD4C,
    16'h4DE4,
    16'h0935,
    16'hAD1A,
    16'hD51C,
    16'h37E8,
    16'hD89B,
    16'h133B,
    16'h4F92,
    16'h7956,
    16'hF200,
    16'h58C5,
    16'h8902,
    16'h301A,
    16'hA87B,
    16'h42F8,
    16'h8CE8,
    16'hD960,
    16'h947C,
    16'h681B,
    16'h5163,
    16'hE2F4,
    16'hA437,
    16'h9D46,
    16'h45BD,
    16'h7D75,
    16'h2313,
    16'h6161,
    16'hBAE4,
    16'h037D,
    16'h9F47,
    16'h1157,
    16'h79F4,
    16'h9059,
    16'h49C9,
    16'hD632,
    16'h23DA,
    16'h536A,
    16'h0A09,
    16'h981F,
    16'h5E85,
    16'h14B8,
    16'h4CEA,
    16'hDDB6,
    16'hAC4E,
    16'h6FEA,
    16'h20B5,
    16'h90D7,
    16'h2665,
    16'h7702,
    16'h9C64,
    16'h9D41,
    16'hC2EA,
    16'h181D,
    16'h797D,
    16'hC98C,
    16'h2951,
    16'hA2FD,
    16'h931D,
    16'h066E,
    16'h451D,
    16'h0760,
    16'h0B9A,
    16'h8AA4,
    16'h69D8,
    16'h8EF7,
    16'h4907,
    16'h3417,
    16'hF905,
    16'h799B,
    16'h17FE,
    16'h1DAA,
    16'h2215,
    16'hA75C,
    16'h1DCA,
    16'h7F33,
    16'h2DDC,
    16'h1015,
    16'hC11E,
    16'hDDD2,
    16'hA437,
    16'h03F1,
    16'h1E1B,
    16'h8765,
    16'h3019,
    16'h50BE,
    16'h1C34,
    16'h5668,
    16'h60D8,
    16'h746A,
    16'h2C8C,
    16'hF295,
    16'h76FD,
    16'hB134,
    16'h2FD5,
    16'hB2E6,
    16'hC941,
    16'h5D35,
    16'h8185,
    16'h4ED0,
    16'h0767,
    16'h31F3,
    16'h4B68,
    16'h9757,
    16'h908E,
    16'h43AC,
    16'h6765,
    16'h494A,
    16'hC448,
    16'h66A2,
    16'h48BF,
    16'h4FA9,
    16'h1FFF,
    16'h9C43,
    16'hFC16,
    16'hDDEA,
    16'hBA93,
    16'h5E9E,
    16'h6102,
    16'h7F2A,
    16'h9E25,
    16'hB4F5,
    16'hC545,
    16'hD089,
    16'hB07D,
    16'h0753,
    16'h0AE6,
    16'h7B4A,
    16'h7FD7,
    16'h48EA,
    16'hEAE6,
    16'h0389,
    16'h23C5,
    16'hFE3E,
    16'h91DB,
    16'h7E95,
    16'h7E56,
    16'h34E8,
    16'h6E95,
    16'hD838,
    16'hB63A,
    16'hADA9,
    16'h23C0,
    16'hA6A9,
    16'hC88E,
    16'h5D37,
    16'hB744,
    16'h4BB3,
    16'h242F,
    16'hF4F4,
    16'h56D4,
    16'hE878,
    16'hDA34,
    16'hE1D0,
    16'h78BE,
    16'hA563,
    16'h6F3C,
    16'h2EC4,
    16'h09AE,
    16'h4FEF,
    16'hFE51,
    16'hA579,
    16'h46A4,
    16'h9175,
    16'hE2A3,
    16'h8847,
    16'h8B9F,
    16'h95FC,
    16'hE9EE,
    16'hB1CD,
    16'h3561,
    16'hBFE9,
    16'hA029,
    16'h4ED1,
    16'h33BE,
    16'h353A,
    16'h47B4,
    16'h3ED6,
    16'h8167,
    16'hAC9F,
    16'h36B4,
    16'h9AD1,
    16'hB445,
    16'h61C8,
    16'hC19F,
    16'h6C3E,
    16'h66C1,
    16'h77DC,
    16'hC466,
    16'h4773,
    16'hB4A7,
    16'h7FC4,
    16'h1ECF,
    16'hB34A,
    16'h5C39,
    16'h4FE7,
    16'h9EFD,
    16'hF1C7,
    16'hF424,
    16'h58AC,
    16'h1A8D,
    16'hA113,
    16'hBAB8,
    16'hCEF1,
    16'h08B5,
    16'h62B0,
    16'hEA76,
    16'hDA8A,
    16'hFA2D,
    16'h5194,
    16'h6C61,
    16'hF0AE,
    16'hB453,
    16'h3407,
    16'h1BD8,
    16'h8581,
    16'h4C20,
    16'hA324,
    16'hF7C8,
    16'hE805,
    16'h0651,
    16'h84AC,
    16'hF1D8,
    16'hA389,
    16'hC2B1,
    16'h4B64,
    16'h5E69,
    16'h62B6,
    16'h989C,
    16'h5B38,
    16'hEBD4,
    16'h6209,
    16'h9721,
    16'hEA24,
    16'h15B5,
    16'h664B,
    16'h327E,
    16'h1141,
    16'hB35B,
    16'hE3D8,
    16'h1122,
    16'h7818,
    16'hD8F3,
    16'h7B14,
    16'hBF79,
    16'hA648,
    16'hE213,
    16'h0FD2,
    16'hEB38,
    16'h4703,
    16'h3E0A,
    16'h90E4,
    16'h4604,
    16'hF7E3,
    16'h1DE8,
    16'hD71E,
    16'hA803,
    16'h7711,
    16'h8B00,
    16'h9D79,
    16'hA677,
    16'hE64A,
    16'h8B39,
    16'h8469,
    16'h3622,
    16'h0480,
    16'h95BC,
    16'hF031,
    16'h00F7,
    16'h58E5,
    16'h370D,
    16'hA251,
    16'h1019,
    16'h7409,
    16'h9941,
    16'hCB71,
    16'h17B3,
    16'h4319,
    16'h1E13
};
bit [15:0] ave_data_rom[0:1023] = {
    16'h0061,
    16'h00D7,
    16'h01E2,
    16'h02A9,
    16'h035B,
    16'h047D,
    16'h05BC,
    16'h05C1,
    16'h06A5,
    16'h07F0,
    16'h08C0,
    16'h09D9,
    16'h0B47,
    16'h0BC9,
    16'h0C49,
    16'h0E02,
    16'h0F18,
    16'h1040,
    16'h1214,
    16'h13B8,
    16'h1442,
    16'h15BB,
    16'h170F,
    16'h18BC,
    16'h18FE,
    16'h1A30,
    16'h1C2C,
    16'h1C96,
    16'h1E1F,
    16'h1E3F,
    16'h1F93,
    16'h1FA2,
    16'h1FA4,
    16'h20BA,
    16'h218C,
    16'h21A2,
    16'h22A0,
    16'h237C,
    16'h24AB,
    16'h256C,
    16'h259B,
    16'h262F,
    16'h2783,
    16'h27B4,
    16'h2836,
    16'h28A7,
    16'h2A28,
    16'h2B9B,
    16'h2CFB,
    16'h2D51,
    16'h2E9B,
    16'h2EBA,
    16'h2FB5,
    16'h30AA,
    16'h30D2,
    16'h31BB,
    16'h31C6,
    16'h31E4,
    16'h31EA,
    16'h3371,
    16'h3383,
    16'h3432,
    16'h34CA,
    16'h3599,
    16'h372C,
    16'h38C6,
    16'h39BD,
    16'h3A17,
    16'h3A82,
    16'h3C61,
    16'h3E1D,
    16'h3E75,
    16'h3FFE,
    16'h41A7,
    16'h4269,
    16'h427E,
    16'h4359,
    16'h448D,
    16'h45EA,
    16'h46F1,
    16'h4853,
    16'h491F,
    16'h49C3,
    16'h49F2,
    16'h4B2B,
    16'h4C50,
    16'h4D1C,
    16'h4D43,
    16'h4E15,
    16'h4F8A,
    16'h5121,
    16'h51CB,
    16'h5394,
    16'h5527,
    16'h552F,
    16'h56DB,
    16'h5893,
    16'h5982,
    16'h5B2B,
    16'h5C43,
    16'h5DDD,
    16'h5EA6,
    16'h5F9F,
    16'h6079,
    16'h6080,
    16'h6179,
    16'h6185,
    16'h6242,
    16'h6245,
    16'h63D3,
    16'h644A,
    16'h6468,
    16'h6644,
    16'h676C,
    16'h680E,
    16'h6951,
    16'h6993,
    16'h6996,
    16'h6A8F,
    16'h6C7E,
    16'h6D65,
    16'h6DE1,
    16'h6E9A,
    16'h6FB7,
    16'h7068,
    16'h714D,
    16'h718F,
    16'h7379,
    16'h73BD,
    16'h73B2,
    16'h7426,
    16'h73D3,
    16'h73E5,
    16'h72FA,
    16'h7225,
    16'h73D8,
    16'h7332,
    16'h73A4,
    16'h7406,
    16'h73DC,
    16'h741A,
    16'h74E0,
    16'h7528,
    16'h73F0,
    16'h73A0,
    16'h7315,
    16'h732C,
    16'h71A6,
    16'h7204,
    16'h714B,
    16'h7087,
    16'h6FC3,
    16'h714F,
    16'h7113,
    16'h6F5C,
    16'h6F1E,
    16'h6F28,
    16'h6F65,
    16'h6FF4,
    16'h703B,
    16'h71AB,
    16'h7185,
    16'h71D2,
    16'h71C8,
    16'h714F,
    16'h721A,
    16'h729A,
    16'h71DB,
    16'h71CC,
    16'h71BF,
    16'h7078,
    16'h7210,
    16'h7205,
    16'h735B,
    16'h734D,
    16'h73BF,
    16'h726D,
    16'h73DC,
    16'h7436,
    16'h75D8,
    16'h7547,
    16'h75F4,
    16'h76D2,
    16'h77A9,
    16'h793E,
    16'h7A1E,
    16'h7BB6,
    16'h7B19,
    16'h7C7A,
    16'h7CF8,
    16'h7CEE,
    16'h7DD9,
    16'h7CF1,
    16'h7C9D,
    16'h7D95,
    16'h7ED6,
    16'h801D,
    16'h7E62,
    16'h7DAE,
    16'h7ECC,
    16'h7D81,
    16'h7C06,
    16'h7D23,
    16'h7D89,
    16'h7E09,
    16'h7DED,
    16'h7D95,
    16'h7E64,
    16'h7E6B,
    16'h7F10,
    16'h7EEB,
    16'h7F05,
    16'h7EFB,
    16'h7E72,
    16'h7F8E,
    16'h7F7E,
    16'h7F36,
    16'h7EB4,
    16'h7D8A,
    16'h7DA8,
    16'h7D0D,
    16'h7CFD,
    16'h7E40,
    16'h7D63,
    16'h7C25,
    16'h7C46,
    16'h7BEE,
    16'h7B81,
    16'h7B34,
    16'h7ACD,
    16'h7B32,
    16'h7BF3,
    16'h7DB3,
    16'h7E61,
    16'h8037,
    16'h8154,
    16'h82FA,
    16'h82C4,
    16'h8325,
    16'h8402,
    16'h831F,
    16'h8301,
    16'h840D,
    16'h8458,
    16'h84EC,
    16'h866E,
    16'h8721,
    16'h864B,
    16'h856A,
    16'h85BF,
    16'h865C,
    16'h86D5,
    16'h879C,
    16'h87E2,
    16'h888D,
    16'h87FE,
    16'h8833,
    16'h891B,
    16'h87D4,
    16'h8913,
    16'h88B7,
    16'h888F,
    16'h890A,
    16'h88B2,
    16'h891F,
    16'h887F,
    16'h88C4,
    16'h87DC,
    16'h8764,
    16'h871E,
    16'h8764,
    16'h87BC,
    16'h88DD,
    16'h8867,
    16'h8792,
    16'h87AF,
    16'h883C,
    16'h8950,
    16'h8955,
    16'h8A42,
    16'h890F,
    16'h887B,
    16'h8924,
    16'h89C7,
    16'h89B7,
    16'h89DD,
    16'h89ED,
    16'h89FF,
    16'h8951,
    16'h8884,
    16'h8855,
    16'h889F,
    16'h8911,
    16'h8962,
    16'h8885,
    16'h8918,
    16'h893E,
    16'h8A3A,
    16'h8A35,
    16'h89B4,
    16'h8A47,
    16'h892F,
    16'h8945,
    16'h88D8,
    16'h88F9,
    16'h88C4,
    16'h8897,
    16'h881E,
    16'h89B4,
    16'h8961,
    16'h88F7,
    16'h88BA,
    16'h8748,
    16'h8711,
    16'h86DF,
    16'h872E,
    16'h8699,
    16'h863E,
    16'h86E4,
    16'h85ED,
    16'h8640,
    16'h859F,
    16'h8482,
    16'h83AF,
    16'h824E,
    16'h837B,
    16'h8390,
    16'h8273,
    16'h82AC,
    16'h8403,
    16'h8337,
    16'h8332,
    16'h82FC,
    16'h83AC,
    16'h82F0,
    16'h8215,
    16'h8183,
    16'h8069,
    16'h8080,
    16'h816C,
    16'h8168,
    16'h8298,
    16'h827F,
    16'h834F,
    16'h835F,
    16'h841B,
    16'h8592,
    16'h8561,
    16'h8484,
    16'h841B,
    16'h8353,
    16'h836F,
    16'h84ED,
    16'h84EC,
    16'h8586,
    16'h84FC,
    16'h851B,
    16'h84D2,
    16'h8517,
    16'h83C4,
    16'h826B,
    16'h82B5,
    16'h81A0,
    16'h8141,
    16'h802C,
    16'h808D,
    16'h819E,
    16'h8132,
    16'h81D9,
    16'h81AE,
    16'h8080,
    16'h8025,
    16'h7F8B,
    16'h7FF4,
    16'h7F7A,
    16'h7FE2,
    16'h819D,
    16'h81B5,
    16'h81C9,
    16'h81CE,
    16'h8144,
    16'h80BB,
    16'h815B,
    16'h80EC,
    16'h813E,
    16'h814C,
    16'h82E9,
    16'h81AA,
    16'h8143,
    16'h825F,
    16'h8214,
    16'h8218,
    16'h81DC,
    16'h829E,
    16'h81DC,
    16'h8284,
    16'h8335,
    16'h833B,
    16'h82A8,
    16'h833B,
    16'h8290,
    16'h8397,
    16'h83E3,
    16'h845B,
    16'h8395,
    16'h837F,
    16'h8480,
    16'h845B,
    16'h8526,
    16'h859C,
    16'h8650,
    16'h868C,
    16'h8579,
    16'h84F5,
    16'h83E9,
    16'h853D,
    16'h84DE,
    16'h85CB,
    16'h8513,
    16'h859A,
    16'h85F0,
    16'h8545,
    16'h84FF,
    16'h8513,
    16'h8656,
    16'h858E,
    16'h86B2,
    16'h8714,
    16'h86C1,
    16'h86E8,
    16'h8650,
    16'h84F7,
    16'h8675,
    16'h85EC,
    16'h84B9,
    16'h83A0,
    16'h8373,
    16'h82EB,
    16'h82D8,
    16'h8228,
    16'h83C7,
    16'h843D,
    16'h839E,
    16'h83CB,
    16'h8340,
    16'h8449,
    16'h848E,
    16'h8497,
    16'h83C4,
    16'h8481,
    16'h851B,
    16'h849A,
    16'h85EC,
    16'h85EA,
    16'h8581,
    16'h85C8,
    16'h85D5,
    16'h857F,
    16'h8587,
    16'h8638,
    16'h8598,
    16'h842D,
    16'h85AB,
    16'h8532,
    16'h852A,
    16'h86A5,
    16'h871D,
    16'h86DC,
    16'h8791,
    16'h867F,
    16'h85F1,
    16'h8668,
    16'h8785,
    16'h876F,
    16'h85A1,
    16'h85E9,
    16'h870E,
    16'h8695,
    16'h878A,
    16'h8749,
    16'h8747,
    16'h87DE,
    16'h862F,
    16'h87F0,
    16'h8851,
    16'h88A3,
    16'h87B0,
    16'h889A,
    16'h8903,
    16'h888F,
    16'h893F,
    16'h89BF,
    16'h89ED,
    16'h89C3,
    16'h8840,
    16'h87DB,
    16'h8804,
    16'h88EE,
    16'h88AA,
    16'h87A9,
    16'h88EC,
    16'h88A7,
    16'h8948,
    16'h88A5,
    16'h8755,
    16'h8796,
    16'h874B,
    16'h8653,
    16'h8579,
    16'h85C4,
    16'h847B,
    16'h83BF,
    16'h83AB,
    16'h83BB,
    16'h821A,
    16'h8239,
    16'h8242,
    16'h814D,
    16'h80C5,
    16'h7FD5,
    16'h80CE,
    16'h7F8C,
    16'h7F88,
    16'h8074,
    16'h7FC6,
    16'h800D,
    16'h80DD,
    16'h80E4,
    16'h8115,
    16'h81A5,
    16'h80C3,
    16'h8158,
    16'h8216,
    16'h805C,
    16'h7FD0,
    16'h7EE1,
    16'h7EF9,
    16'h7E6B,
    16'h7D51,
    16'h7DC4,
    16'h7D7E,
    16'h7E2E,
    16'h7E9E,
    16'h7EA9,
    16'h7F80,
    16'h8037,
    16'h81FB,
    16'h81EC,
    16'h8264,
    16'h8122,
    16'h824A,
    16'h833E,
    16'h82A0,
    16'h833F,
    16'h83B9,
    16'h8350,
    16'h8405,
    16'h8524,
    16'h8612,
    16'h87DD,
    16'h8689,
    16'h858A,
    16'h85F8,
    16'h8788,
    16'h87AD,
    16'h877F,
    16'h8700,
    16'h87FD,
    16'h8801,
    16'h8724,
    16'h8796,
    16'h86A0,
    16'h8816,
    16'h8828,
    16'h8822,
    16'h892D,
    16'h8A38,
    16'h8A25,
    16'h8990,
    16'h8B14,
    16'h8991,
    16'h8A09,
    16'h8AD4,
    16'h8A7A,
    16'h8A77,
    16'h8A07,
    16'h89EC,
    16'h8A40,
    16'h8A25,
    16'h8BC4,
    16'h8A5B,
    16'h8BA1,
    16'h8ADE,
    16'h8A75,
    16'h8B3C,
    16'h8B9C,
    16'h8B09,
    16'h8C14,
    16'h8C3E,
    16'h8BD6,
    16'h8A31,
    16'h89D8,
    16'h8AD6,
    16'h8AEF,
    16'h8AED,
    16'h8B46,
    16'h8A5C,
    16'h8AAF,
    16'h8A32,
    16'h897F,
    16'h8ACE,
    16'h8918,
    16'h8759,
    16'h8720,
    16'h8748,
    16'h8637,
    16'h85FC,
    16'h861F,
    16'h852A,
    16'h8428,
    16'h850E,
    16'h841C,
    16'h83F7,
    16'h84D8,
    16'h84B0,
    16'h8324,
    16'h832C,
    16'h8311,
    16'h8344,
    16'h82C8,
    16'h8147,
    16'h8136,
    16'h8271,
    16'h81D8,
    16'h824D,
    16'h82C7,
    16'h83A3,
    16'h847E,
    16'h8484,
    16'h85CA,
    16'h8549,
    16'h8593,
    16'h85AA,
    16'h85BF,
    16'h8766,
    16'h8853,
    16'h89DB,
    16'h8B29,
    16'h8A7E,
    16'h8AAD,
    16'h8B21,
    16'h8A89,
    16'h8AC8,
    16'h8A1F,
    16'h8AA7,
    16'h8AE3,
    16'h89C1,
    16'h89DA,
    16'h8B21,
    16'h8AD2,
    16'h8A88,
    16'h8BC2,
    16'h8BB4,
    16'h8C6A,
    16'h8B8A,
    16'h8B8F,
    16'h8B64,
    16'h8A87,
    16'h8B33,
    16'h8B18,
    16'h8B55,
    16'h8A38,
    16'h89CC,
    16'h89E8,
    16'h890B,
    16'h88DE,
    16'h8902,
    16'h8982,
    16'h87EF,
    16'h880D,
    16'h891A,
    16'h8997,
    16'h8949,
    16'h8825,
    16'h86C8,
    16'h8562,
    16'h8426,
    16'h833A,
    16'h849C,
    16'h85CE,
    16'h864E,
    16'h8519,
    16'h84E7,
    16'h856D,
    16'h862C,
    16'h8546,
    16'h83AE,
    16'h8513,
    16'h85C3,
    16'h873A,
    16'h8692,
    16'h8676,
    16'h85C7,
    16'h844D,
    16'h844C,
    16'h84F3,
    16'h846D,
    16'h8448,
    16'h844C,
    16'h82B5,
    16'h8290,
    16'h834B,
    16'h843A,
    16'h8433,
    16'h8362,
    16'h82E4,
    16'h82D6,
    16'h81CA,
    16'h81DF,
    16'h801B,
    16'h8051,
    16'h7FF1,
    16'h7E44,
    16'h7EEC,
    16'h7EE3,
    16'h7E75,
    16'h7D21,
    16'h7CD8,
    16'h7DCF,
    16'h7DFB,
    16'h7D5E,
    16'h7D97,
    16'h7DDF,
    16'h7DAD,
    16'h7EDF,
    16'h7E0F,
    16'h7CFD,
    16'h7D47,
    16'h7C37,
    16'h7CD5,
    16'h7E91,
    16'h7FA9,
    16'h7F53,
    16'h7F96,
    16'h8071,
    16'h80CB,
    16'h80DE,
    16'h7FF6,
    16'h7FAB,
    16'h80B6,
    16'h80E6,
    16'h818C,
    16'h8011,
    16'h8074,
    16'h8122,
    16'h82F0,
    16'h81EF,
    16'h81D3,
    16'h81E2,
    16'h8267,
    16'h8140,
    16'h81C9,
    16'h81E7,
    16'h81F3,
    16'h81D5,
    16'h80AF,
    16'h822C,
    16'h81FD,
    16'h829E,
    16'h8171,
    16'h8220,
    16'h81BF,
    16'h80D0,
    16'h8123,
    16'h7F90,
    16'h7F0D,
    16'h7E73,
    16'h7E9B,
    16'h7E96,
    16'h7E26,
    16'h7E5D,
    16'h7DFE,
    16'h7CD2,
    16'h7B38,
    16'h7C1C,
    16'h7B03,
    16'h7966,
    16'h7906,
    16'h799D,
    16'h79B8,
    16'h799D,
    16'h7867,
    16'h78EA,
    16'h78E7,
    16'h7979,
    16'h7A11,
    16'h7A76,
    16'h7B66,
    16'h7A04,
    16'h7A4C,
    16'h7B0F,
    16'h797F,
    16'h79A5,
    16'h7A2B,
    16'h7850,
    16'h784F,
    16'h783D,
    16'h7699,
    16'h75B6,
    16'h74B2,
    16'h7478,
    16'h74ED,
    16'h7547,
    16'h76A9,
    16'h76FA,
    16'h762C,
    16'h74AC,
    16'h73B5,
    16'h73D2,
    16'h7384,
    16'h72BC,
    16'h71FB,
    16'h714F,
    16'h71EA,
    16'h736B,
    16'h72EF,
    16'h7108,
    16'h6F5D,
    16'h6F4B,
    16'h6DDA,
    16'h6DB8,
    16'h6D92,
    16'h6D0C,
    16'h6BD5,
    16'h6C6E,
    16'h6B23,
    16'h6CE2,
    16'h6DA1,
    16'h6DA9,
    16'h6D08,
    16'h6CFD,
    16'h6DD7,
    16'h6E62,
    16'h6E69,
    16'h6EAB,
    16'h6DC9,
    16'h6DBA,
    16'h6E4E,
    16'h6F3A,
    16'h6F51,
    16'h6FB2,
    16'h6E85,
    16'h6DD2,
    16'h6E03,
    16'h6EBA,
    16'h6E9F,
    16'h6E35,
    16'h6D0A,
    16'h6DCB,
    16'h6E93,
    16'h6E92,
    16'h6F41,
    16'h6E3C,
    16'h6ED0,
    16'h6F69,
    16'h6F67,
    16'h7056,
    16'h7117,
    16'h70F0,
    16'h7105,
    16'h7092,
    16'h7045,
    16'h6FC5,
    16'h6ECA,
    16'h6EC0,
    16'h7083,
    16'h6F30,
    16'h6DCD,
    16'h6F5A,
    16'h6ECC,
    16'h6FA3,
    16'h7001,
    16'h6F78,
    16'h6E71,
    16'h6F70,
    16'h6FCA,
    16'h70C5,
    16'h6FBC,
    16'h7083,
    16'h70FB,
    16'h7002,
    16'h7048,
    16'h700F,
    16'h6FB5,
    16'h6FD9,
    16'h6F3E,
    16'h6FD4,
    16'h70FD,
    16'h71C6,
    16'h7271,
    16'h72F9,
    16'h7262,
    16'h72B9,
    16'h718D,
    16'h720B,
    16'h7313,
    16'h733D,
    16'h7337,
    16'h72AE,
    16'h742B,
    16'h7495,
    16'h7598,
    16'h7594,
    16'h76AB,
    16'h77E5,
    16'h77B6,
    16'h777A,
    16'h7762,
    16'h7720,
    16'h7746,
    16'h768F,
    16'h76D1,
    16'h7661,
    16'h762B,
    16'h764A,
    16'h7531,
    16'h7637,
    16'h76AC,
    16'h75DD,
    16'h770D,
    16'h76A0,
    16'h7647,
    16'h772A,
    16'h7828,
    16'h78A9,
    16'h79FB,
    16'h79E5,
    16'h794F,
    16'h7998,
    16'h79BE,
    16'h79F6,
    16'h7941,
    16'h7A32,
    16'h7BEA,
    16'h7C60,
    16'h7C51,
    16'h7C45,
    16'h7D7E,
    16'h7E1E,
    16'h7DD4,
    16'h7E79,
    16'h7ECB,
    16'h7EC5,
    16'h7F71,
    16'h800C,
    16'h80A9,
    16'h817B,
    16'h8284,
    16'h824A,
    16'h824A,
    16'h82A8,
    16'h827E,
    16'h82DC,
    16'h8472,
    16'h845D,
    16'h837C,
    16'h8323,
    16'h84A7,
    16'h8488,
    16'h847B,
    16'h8457,
    16'h8411,
    16'h8439,
    16'h855B,
    16'h85AE,
    16'h86EF,
    16'h8684,
    16'h8691,
    16'h87DE,
    16'h873B,
    16'h8775,
    16'h8651,
    16'h85A6,
    16'h867C,
    16'h87A4,
    16'h8786,
    16'h873E,
    16'h86F8,
    16'h8632,
    16'h863C,
    16'h86CB,
    16'h87CD,
    16'h86EE,
    16'h8789,
    16'h86AD,
    16'h859E,
    16'h851F,
    16'h844A,
    16'h862B,
    16'h8651,
    16'h8709,
    16'h8759,
    16'h87B5,
    16'h86F6,
    16'h882A,
    16'h892F,
    16'h88FF,
    16'h88F2,
    16'h88FD,
    16'h886D,
    16'h880C,
    16'h885B,
    16'h888A,
    16'h8720,
    16'h8676,
    16'h869D,
    16'h8694,
    16'h8523,
    16'h8551,
    16'h8515,
    16'h8615,
    16'h85FC,
    16'h8498,
    16'h8426
};

int raw_file;
int ave_file;
string raw_line;
string ave_line;
int raw_count = 1;
int ave_count = 1;

// module
MOVING_AVE U_MOVING_AVE(
.*,
.ASI_READY(ASI_READY),
.ASI_VALID(ASI_VALID),
.ASI_DATA(ASI_DATA),
.ASO_VALID(ASO_VALID),
.ASO_DATA(ASO_DATA),
.ASO_ERROR(ASO_ERROR)
);


/*=============================================================================
 * Clock
 *============================================================================*/
always begin
    #(ClkCyc);
    CLK = ~CLK;
end


/*=============================================================================
 * Reset
 *============================================================================*/
initial begin
    #(ResetTime);
    RESET_n = 1;
end 


/*=============================================================================
 * Signal initialization
 *============================================================================*/
initial begin
    ASI_VALID = 1'b0;
    ASI_DATA = 16'd0;

    #(ResetTime);
    @(posedge CLK);

/*=============================================================================
 * Data check
 *============================================================================*/
    $display("%0s(%0d)Normalized data check", `__FILE__, `__LINE__);
    wait(ASI_READY);
    ASI_DATA = 0;
    @(posedge CLK);
    ASI_VALID = 1'b1;
    for (int i=0;i<128;i++) begin
        ASI_DATA = 16'h7fff;
        @(posedge CLK);
    end
    for (int i=0;i<18;i++) begin
        @(posedge CLK);
    end

    @(posedge CLK);
    ASI_DATA = 0;
    ASI_VALID = 1'b0;
    @(posedge CLK);
    RESET_n = 0;
    @(posedge CLK);
    RESET_n = 1;

    $display("%0s(%0d)Normal data check", `__FILE__, `__LINE__);
    wait(ASI_READY);
    @(posedge CLK);
    ASI_VALID = 1'b1;
    for (int i=0;i<1024;i++) begin
        ASI_DATA = raw_data_rom[i];
        @(posedge CLK);
    end
end

initial begin
    wait(ASO_VALID);
    for (int i=0;i<128;i++) begin
        @(posedge CLK);
    end
    for (int i=0;i<10;i++) begin
        wait(ASO_VALID);
        @(negedge CLK);
        `ChkValue("ASO_DATA", ASO_DATA, 16'h7fff);
    end
    for (int i=0;i<10;i++) begin
        @(posedge CLK);
    end
    for (int i=0;i<1024;i++) begin
        wait(ASO_VALID);
        @(negedge CLK);
        `ChkValue("ASO_DATA", ASO_DATA, ave_data_rom[i]);
    end

    $finish;
end

endmodule
// TB_MOVING_AVE